`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    12:34:59 11/28/2017 
// Design Name: 
// Module Name:    divisions_lut 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module divisions_lut(
    input [8:0] M,
    output reg [16:0] out
    );

	always @ * begin
		case (M)
					9'b000000001: out = 16'b1111111111111111;
					9'b000000010: out = 16'b0111111111111111;
					9'b000000011: out = 16'b0101010101010101;
					9'b000000100: out = 16'b0011111111111111;
					9'b000000101: out = 16'b0011001100110011;
					9'b000000110: out = 16'b0010101010101010;
					9'b000000111: out = 16'b0010010010010010;
					9'b000001000: out = 16'b0001111111111111;
					9'b000001001: out = 16'b0001110001110001;
					9'b000001010: out = 16'b0001100110011001;
					9'b000001011: out = 16'b0001011101000101;
					9'b000001100: out = 16'b0001010101010101;
					9'b000001101: out = 16'b0001001110110001;
					9'b000001110: out = 16'b0001001001001001;
					9'b000001111: out = 16'b0001000100010001;
					9'b000010000: out = 16'b0000111111111111;
					9'b000010001: out = 16'b0000111100001111;
					9'b000010010: out = 16'b0000111000111000;
					9'b000010011: out = 16'b0000110101111001;
					9'b000010100: out = 16'b0000110011001100;
					9'b000010101: out = 16'b0000110000110000;
					9'b000010110: out = 16'b0000101110100010;
					9'b000010111: out = 16'b0000101100100001;
					9'b000011000: out = 16'b0000101010101010;
					9'b000011001: out = 16'b0000101000111101;
					9'b000011010: out = 16'b0000100111011000;
					9'b000011011: out = 16'b0000100101111011;
					9'b000011100: out = 16'b0000100100100100;
					9'b000011101: out = 16'b0000100011010011;
					9'b000011110: out = 16'b0000100010001000;
					9'b000011111: out = 16'b0000100001000010;
					9'b000100000: out = 16'b0000011111111111;
					9'b000100001: out = 16'b0000011111000001;
					9'b000100010: out = 16'b0000011110000111;
					9'b000100011: out = 16'b0000011101010000;
					9'b000100100: out = 16'b0000011100011100;
					9'b000100101: out = 16'b0000011011101011;
					9'b000100110: out = 16'b0000011010111100;
					9'b000100111: out = 16'b0000011010010000;
					9'b000101000: out = 16'b0000011001100110;
					9'b000101001: out = 16'b0000011000111110;
					9'b000101010: out = 16'b0000011000011000;
					9'b000101011: out = 16'b0000010111110100;
					9'b000101100: out = 16'b0000010111010001;
					9'b000101101: out = 16'b0000010110110000;
					9'b000101110: out = 16'b0000010110010000;
					9'b000101111: out = 16'b0000010101110010;
					9'b000110000: out = 16'b0000010101010101;
					9'b000110001: out = 16'b0000010100111001;
					9'b000110010: out = 16'b0000010100011110;
					9'b000110011: out = 16'b0000010100000101;
					9'b000110100: out = 16'b0000010011101100;
					9'b000110101: out = 16'b0000010011010100;
					9'b000110110: out = 16'b0000010010111101;
					9'b000110111: out = 16'b0000010010100111;
					9'b000111000: out = 16'b0000010010010010;
					9'b000111001: out = 16'b0000010001111101;
					9'b000111010: out = 16'b0000010001101001;
					9'b000111011: out = 16'b0000010001010110;
					9'b000111100: out = 16'b0000010001000100;
					9'b000111101: out = 16'b0000010000110010;
					9'b000111110: out = 16'b0000010000100001;
					9'b000111111: out = 16'b0000010000010000;
					9'b001000000: out = 16'b0000001111111111;
					9'b001000001: out = 16'b0000001111110000;
					9'b001000010: out = 16'b0000001111100000;
					9'b001000011: out = 16'b0000001111010010;
					9'b001000100: out = 16'b0000001111000011;
					9'b001000101: out = 16'b0000001110110101;
					9'b001000110: out = 16'b0000001110101000;
					9'b001000111: out = 16'b0000001110011011;
					9'b001001000: out = 16'b0000001110001110;
					9'b001001001: out = 16'b0000001110000001;
					9'b001001010: out = 16'b0000001101110101;
					9'b001001011: out = 16'b0000001101101001;
					9'b001001100: out = 16'b0000001101011110;
					9'b001001101: out = 16'b0000001101010011;
					9'b001001110: out = 16'b0000001101001000;
					9'b001001111: out = 16'b0000001100111101;
					9'b001010000: out = 16'b0000001100110011;
					9'b001010001: out = 16'b0000001100101001;
					9'b001010010: out = 16'b0000001100011111;
					9'b001010011: out = 16'b0000001100010101;
					9'b001010100: out = 16'b0000001100001100;
					9'b001010101: out = 16'b0000001100000011;
					9'b001010110: out = 16'b0000001011111010;
					9'b001010111: out = 16'b0000001011110001;
					9'b001011000: out = 16'b0000001011101000;
					9'b001011001: out = 16'b0000001011100000;
					9'b001011010: out = 16'b0000001011011000;
					9'b001011011: out = 16'b0000001011010000;
					9'b001011100: out = 16'b0000001011001000;
					9'b001011101: out = 16'b0000001011000000;
					9'b001011110: out = 16'b0000001010111001;
					9'b001011111: out = 16'b0000001010110001;
					9'b001100000: out = 16'b0000001010101010;
					9'b001100001: out = 16'b0000001010100011;
					9'b001100010: out = 16'b0000001010011100;
					9'b001100011: out = 16'b0000001010010101;
					9'b001100100: out = 16'b0000001010001111;
					9'b001100101: out = 16'b0000001010001000;
					9'b001100110: out = 16'b0000001010000010;
					9'b001100111: out = 16'b0000001001111100;
					9'b001101000: out = 16'b0000001001110110;
					9'b001101001: out = 16'b0000001001110000;
					9'b001101010: out = 16'b0000001001101010;
					9'b001101011: out = 16'b0000001001100100;
					9'b001101100: out = 16'b0000001001011110;
					9'b001101101: out = 16'b0000001001011001;
					9'b001101110: out = 16'b0000001001010011;
					9'b001101111: out = 16'b0000001001001110;
					9'b001110000: out = 16'b0000001001001001;
					9'b001110001: out = 16'b0000001001000011;
					9'b001110010: out = 16'b0000001000111110;
					9'b001110011: out = 16'b0000001000111001;
					9'b001110100: out = 16'b0000001000110100;
					9'b001110101: out = 16'b0000001000110000;
					9'b001110110: out = 16'b0000001000101011;
					9'b001110111: out = 16'b0000001000100110;
					9'b001111000: out = 16'b0000001000100010;
					9'b001111001: out = 16'b0000001000011101;
					9'b001111010: out = 16'b0000001000011001;
					9'b001111011: out = 16'b0000001000010100;
					9'b001111100: out = 16'b0000001000010000;
					9'b001111101: out = 16'b0000001000001100;
					9'b001111110: out = 16'b0000001000001000;
					9'b001111111: out = 16'b0000001000000100;
					9'b010000000: out = 16'b0000000111111111;
					9'b010000001: out = 16'b0000000111111100;
					9'b010000010: out = 16'b0000000111111000;
					9'b010000011: out = 16'b0000000111110100;
					9'b010000100: out = 16'b0000000111110000;
					9'b010000101: out = 16'b0000000111101100;
					9'b010000110: out = 16'b0000000111101001;
					9'b010000111: out = 16'b0000000111100101;
					9'b010001000: out = 16'b0000000111100001;
					9'b010001001: out = 16'b0000000111011110;
					9'b010001010: out = 16'b0000000111011010;
					9'b010001011: out = 16'b0000000111010111;
					9'b010001100: out = 16'b0000000111010100;
					9'b010001101: out = 16'b0000000111010000;
					9'b010001110: out = 16'b0000000111001101;
					9'b010001111: out = 16'b0000000111001010;
					9'b010010000: out = 16'b0000000111000111;
					9'b010010001: out = 16'b0000000111000011;
					9'b010010010: out = 16'b0000000111000000;
					9'b010010011: out = 16'b0000000110111101;
					9'b010010100: out = 16'b0000000110111010;
					9'b010010101: out = 16'b0000000110110111;
					9'b010010110: out = 16'b0000000110110100;
					9'b010010111: out = 16'b0000000110110010;
					9'b010011000: out = 16'b0000000110101111;
					9'b010011001: out = 16'b0000000110101100;
					9'b010011010: out = 16'b0000000110101001;
					9'b010011011: out = 16'b0000000110100110;
					9'b010011100: out = 16'b0000000110100100;
					9'b010011101: out = 16'b0000000110100001;
					9'b010011110: out = 16'b0000000110011110;
					9'b010011111: out = 16'b0000000110011100;
					9'b010100000: out = 16'b0000000110011001;
					9'b010100001: out = 16'b0000000110010111;
					9'b010100010: out = 16'b0000000110010100;
					9'b010100011: out = 16'b0000000110010010;
					9'b010100100: out = 16'b0000000110001111;
					9'b010100101: out = 16'b0000000110001101;
					9'b010100110: out = 16'b0000000110001010;
					9'b010100111: out = 16'b0000000110001000;
					9'b010101000: out = 16'b0000000110000110;
					9'b010101001: out = 16'b0000000110000011; 
					default: 	  out = 16'b0000000000000000;
		endcase
	end

endmodule
