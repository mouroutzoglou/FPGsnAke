module s_h_d_rom(
        input wire clk,
        input wire [4:0] x,
        input wire [4:0] y,
        output reg [23:0] data
	);
	
	always @ * begin
	case ({y, x})
                10'b0000000000: data = 24'b000000000000000000000000;
                10'b0000000001: data = 24'b000011110000111100001111;
                10'b0000000010: data = 24'b001101010011111100110100;
                10'b0000000011: data = 24'b010111010111111001011011;
                10'b0000000100: data = 24'b010101110111100001010110;
                10'b0000000101: data = 24'b011010001001010001100111;
                10'b0000000110: data = 24'b011101011010011101110011;
                10'b0000000111: data = 24'b011100111010010001110001;
                10'b0000001000: data = 24'b011100111010001101110001;
                10'b0000001001: data = 24'b011101001010011101110010;
                10'b0000001010: data = 24'b011110111011101001111001;
                10'b0000001011: data = 24'b011110111011101001111001;
                10'b0000001100: data = 24'b011110111011101001111001;
                10'b0000001101: data = 24'b011110111011101001111001;
                10'b0000001110: data = 24'b011110111011101001111001;
                10'b0000001111: data = 24'b011110111011101001111001;
                10'b0000010000: data = 24'b011110111011101001111001;
                10'b0000010001: data = 24'b011110111011101001111001;
                10'b0000010010: data = 24'b011110111011101001111001;
                10'b0000010011: data = 24'b011110111011101001111001;
                10'b0000010100: data = 24'b011110111011101001111001;
                10'b0000010101: data = 24'b011110111011101001111001;
                10'b0000010110: data = 24'b011101001010011101110010;
                10'b0000010111: data = 24'b011100111010001101110001;
                10'b0000011000: data = 24'b011100111010010001110001;
                10'b0000011001: data = 24'b011101011010011101110011;
                10'b0000011010: data = 24'b011010001001010001100111;
                10'b0000011011: data = 24'b010101110111100001010110;
                10'b0000011100: data = 24'b010111010111111001011011;
                10'b0000011101: data = 24'b001101010011111100110100;
                10'b0000011110: data = 24'b000011110000111100001111;
                10'b0000011111: data = 24'b000000000000000000000000;
                10'b0000100000: data = 24'b000000000000000000000000;
                10'b0000100001: data = 24'b000000010000000100000001;
                10'b0000100010: data = 24'b001111000101001100111100;
                10'b0000100011: data = 24'b010100000111011001001111;
                10'b0000100100: data = 24'b010011100111001101001101;
                10'b0000100101: data = 24'b011001111001100101100101;
                10'b0000100110: data = 24'b011010101001111101101000;
                10'b0000100111: data = 24'b011010101001111001101000;
                10'b0000101000: data = 24'b011010101001110001101000;
                10'b0000101001: data = 24'b011011011010011101101011;
                10'b0000101010: data = 24'b011101001011011101110010;
                10'b0000101011: data = 24'b011100111011011001110001;
                10'b0000101100: data = 24'b011100111011011001110001;
                10'b0000101101: data = 24'b011100111011011001110001;
                10'b0000101110: data = 24'b011100111011011001110001;
                10'b0000101111: data = 24'b011100111011011001110001;
                10'b0000110000: data = 24'b011100111011011001110001;
                10'b0000110001: data = 24'b011100111011011001110001;
                10'b0000110010: data = 24'b011100111011011001110001;
                10'b0000110011: data = 24'b011100111011011001110001;
                10'b0000110100: data = 24'b011100111011011001110001;
                10'b0000110101: data = 24'b011101001011011101110010;
                10'b0000110110: data = 24'b011011101010100001101100;
                10'b0000110111: data = 24'b011010101001110001101000;
                10'b0000111000: data = 24'b011010101001111001101000;
                10'b0000111001: data = 24'b011010101001111101101000;
                10'b0000111010: data = 24'b011001111001100101100101;
                10'b0000111011: data = 24'b010011100111001101001101;
                10'b0000111100: data = 24'b010100000111011001001111;
                10'b0000111101: data = 24'b001110100101000100111010;
                10'b0000111110: data = 24'b000000000000000000000000;
                10'b0000111111: data = 24'b000000000000000000000000;
                10'b0001000000: data = 24'b000000000000000000000000;
                10'b0001000001: data = 24'b000001100000100000000110;
                10'b0001000010: data = 24'b010011010110111001001101;
                10'b0001000011: data = 24'b010011000110111101001011;
                10'b0001000100: data = 24'b010101100111111101010100;
                10'b0001000101: data = 24'b011010111010000001101001;
                10'b0001000110: data = 24'b011010101001111001101000;
                10'b0001000111: data = 24'b011010101001111001101000;
                10'b0001001000: data = 24'b011010101001110101101000;
                10'b0001001001: data = 24'b011100001010111001101110;
                10'b0001001010: data = 24'b011101001011011101110010;
                10'b0001001011: data = 24'b011100111011011001110001;
                10'b0001001100: data = 24'b011100111011011001110001;
                10'b0001001101: data = 24'b011100111011011001110001;
                10'b0001001110: data = 24'b011100111011011001110001;
                10'b0001001111: data = 24'b011100111011011001110001;
                10'b0001010000: data = 24'b011100111011011001110001;
                10'b0001010001: data = 24'b011100111011011001110001;
                10'b0001010010: data = 24'b011100111011011001110001;
                10'b0001010011: data = 24'b011100111011011001110001;
                10'b0001010100: data = 24'b011100111011011001110001;
                10'b0001010101: data = 24'b011101001011011101110010;
                10'b0001010110: data = 24'b011100001010111001101110;
                10'b0001010111: data = 24'b011010101001110101101000;
                10'b0001011000: data = 24'b011010101001111001101000;
                10'b0001011001: data = 24'b011010101001111001101000;
                10'b0001011010: data = 24'b011010111010000001101001;
                10'b0001011011: data = 24'b010101010111111101010100;
                10'b0001011100: data = 24'b010011000110111101001011;
                10'b0001011101: data = 24'b010011010110111001001101;
                10'b0001011110: data = 24'b000001100000100000000110;
                10'b0001011111: data = 24'b000000000000000000000000;
                10'b0001100000: data = 24'b000000000000000000000000;
                10'b0001100001: data = 24'b001000110010101100100011;
                10'b0001100010: data = 24'b010011110111001001001110;
                10'b0001100011: data = 24'b010011000110111101001011;
                10'b0001100100: data = 24'b010111101000110001011101;
                10'b0001100101: data = 24'b011011001010000101101010;
                10'b0001100110: data = 24'b011010101001111001101000;
                10'b0001100111: data = 24'b011010101001111001101000;
                10'b0001101000: data = 24'b011010101010000001101000;
                10'b0001101001: data = 24'b011100111011010001110001;
                10'b0001101010: data = 24'b011100111011011101110001;
                10'b0001101011: data = 24'b011100111011011001110001;
                10'b0001101100: data = 24'b011100111011011001110001;
                10'b0001101101: data = 24'b011100111011011001110001;
                10'b0001101110: data = 24'b011100111011011001110001;
                10'b0001101111: data = 24'b011100111011011001110001;
                10'b0001110000: data = 24'b011100111011011001110001;
                10'b0001110001: data = 24'b011100111011011001110001;
                10'b0001110010: data = 24'b011100111011011001110001;
                10'b0001110011: data = 24'b011100111011011001110001;
                10'b0001110100: data = 24'b011100111011011001110001;
                10'b0001110101: data = 24'b011100111011011001110001;
                10'b0001110110: data = 24'b011100111011010001110001;
                10'b0001110111: data = 24'b011010101001111101101000;
                10'b0001111000: data = 24'b011010101001111001101000;
                10'b0001111001: data = 24'b011010101001111001101000;
                10'b0001111010: data = 24'b011011001010000101101010;
                10'b0001111011: data = 24'b010111101000110001011101;
                10'b0001111100: data = 24'b010011000110111101001011;
                10'b0001111101: data = 24'b010011110111001001001110;
                10'b0001111110: data = 24'b001001000010101100100100;
                10'b0001111111: data = 24'b000000000000000000000000;
                10'b0010000000: data = 24'b000000000000000000000000;
                10'b0010000001: data = 24'b001011010011110100101101;
                10'b0010000010: data = 24'b010101000111100101010011;
                10'b0010000011: data = 24'b010011000111000101001011;
                10'b0010000100: data = 24'b011001001001010001100010;
                10'b0010000101: data = 24'b011010111001111101101001;
                10'b0010000110: data = 24'b011010101001111001101000;
                10'b0010000111: data = 24'b011010011001110101100111;
                10'b0010001000: data = 24'b011011011010011001101011;
                10'b0010001001: data = 24'b011100111011011101110001;
                10'b0010001010: data = 24'b011100111011011001110001;
                10'b0010001011: data = 24'b011100111011011001110001;
                10'b0010001100: data = 24'b011100111011011001110001;
                10'b0010001101: data = 24'b011100111011011001110001;
                10'b0010001110: data = 24'b011100111011011001110001;
                10'b0010001111: data = 24'b011100111011011001110001;
                10'b0010010000: data = 24'b011100111011011001110001;
                10'b0010010001: data = 24'b011100111011011001110001;
                10'b0010010010: data = 24'b011100111011011001110001;
                10'b0010010011: data = 24'b011100111011011001110001;
                10'b0010010100: data = 24'b011100111011011001110001;
                10'b0010010101: data = 24'b011100111011011001110001;
                10'b0010010110: data = 24'b011100111011011001110001;
                10'b0010010111: data = 24'b011011001010010001101010;
                10'b0010011000: data = 24'b011010101001110101101000;
                10'b0010011001: data = 24'b011010101001111001101000;
                10'b0010011010: data = 24'b011010111001111101101001;
                10'b0010011011: data = 24'b011001001001010001100010;
                10'b0010011100: data = 24'b010011000111000101001011;
                10'b0010011101: data = 24'b010101000111100101010011;
                10'b0010011110: data = 24'b001011000011110000101100;
                10'b0010011111: data = 24'b000000000000000000000000;
                10'b0010100000: data = 24'b000000000000000000000000;
                10'b0010100001: data = 24'b001001110011101000100111;
                10'b0010100010: data = 24'b010100010111100001010000;
                10'b0010100011: data = 24'b010011100111001001001101;
                10'b0010100100: data = 24'b011010001001101001100110;
                10'b0010100101: data = 24'b011010111001111101101001;
                10'b0010100110: data = 24'b011010101001111001101000;
                10'b0010100111: data = 24'b011010011001110101100111;
                10'b0010101000: data = 24'b011100001010110101101110;
                10'b0010101001: data = 24'b011100111011100001110001;
                10'b0010101010: data = 24'b011100111011011001110001;
                10'b0010101011: data = 24'b011100111011011001110001;
                10'b0010101100: data = 24'b011100111011011001110001;
                10'b0010101101: data = 24'b011100111011011001110001;
                10'b0010101110: data = 24'b011100111011011001110001;
                10'b0010101111: data = 24'b011100111011011001110001;
                10'b0010110000: data = 24'b011100111011011001110001;
                10'b0010110001: data = 24'b011100111011011001110001;
                10'b0010110010: data = 24'b011100111011011001110001;
                10'b0010110011: data = 24'b011100111011011001110001;
                10'b0010110100: data = 24'b011100111011011001110001;
                10'b0010110101: data = 24'b011100111011011001110001;
                10'b0010110110: data = 24'b011101001011011101110010;
                10'b0010110111: data = 24'b011011111010101001101101;
                10'b0010111000: data = 24'b011010011001110101100111;
                10'b0010111001: data = 24'b011010101001111001101000;
                10'b0010111010: data = 24'b011010111001111101101001;
                10'b0010111011: data = 24'b011010001001101001100110;
                10'b0010111100: data = 24'b010011100111001001001101;
                10'b0010111101: data = 24'b010100010111100001010000;
                10'b0010111110: data = 24'b001001110011101000100111;
                10'b0010111111: data = 24'b000000000000000000000000;
                10'b0011000000: data = 24'b000000000000000000000000;
                10'b0011000001: data = 24'b001110000100101100111000;
                10'b0011000010: data = 24'b010100000111011001001111;
                10'b0011000011: data = 24'b010100000111011001001111;
                10'b0011000100: data = 24'b011010011001110001100111;
                10'b0011000101: data = 24'b011010101001111101101000;
                10'b0011000110: data = 24'b011010101001111001101000;
                10'b0011000111: data = 24'b011010101001111101101000;
                10'b0011001000: data = 24'b011100101011001101110000;
                10'b0011001001: data = 24'b011100111011011001110001;
                10'b0011001010: data = 24'b011100111011011001110001;
                10'b0011001011: data = 24'b011100111011011001110001;
                10'b0011001100: data = 24'b011100111011011001110001;
                10'b0011001101: data = 24'b011100111011011001110001;
                10'b0011001110: data = 24'b011100111011011001110001;
                10'b0011001111: data = 24'b011100111011011001110001;
                10'b0011010000: data = 24'b011100111011011001110001;
                10'b0011010001: data = 24'b011100111011011001110001;
                10'b0011010010: data = 24'b011100111011011001110001;
                10'b0011010011: data = 24'b011100111011011001110001;
                10'b0011010100: data = 24'b011100111011011001110001;
                10'b0011010101: data = 24'b011100111011011001110001;
                10'b0011010110: data = 24'b011100111011011101110001;
                10'b0011010111: data = 24'b011100011010111101101111;
                10'b0011011000: data = 24'b011010101001110101101000;
                10'b0011011001: data = 24'b011010101001111001101000;
                10'b0011011010: data = 24'b011010101001111101101000;
                10'b0011011011: data = 24'b011010011001110001100111;
                10'b0011011100: data = 24'b010100000111011001001111;
                10'b0011011101: data = 24'b010100000111011001001111;
                10'b0011011110: data = 24'b001110000100101100111000;
                10'b0011011111: data = 24'b000000000000000000000000;
                10'b0011100000: data = 24'b000000000000000000000000;
                10'b0011100001: data = 24'b010001000101101001000100;
                10'b0011100010: data = 24'b010011110111010101001110;
                10'b0011100011: data = 24'b010100010111100001010000;
                10'b0011100100: data = 24'b011010011001110101100111;
                10'b0011100101: data = 24'b011010101001111101101000;
                10'b0011100110: data = 24'b011010101001110101101000;
                10'b0011100111: data = 24'b011011001010001101101010;
                10'b0011101000: data = 24'b011100111011011001110001;
                10'b0011101001: data = 24'b011100111011011001110001;
                10'b0011101010: data = 24'b011100111011011001110001;
                10'b0011101011: data = 24'b011100111011011001110001;
                10'b0011101100: data = 24'b011100111011011001110001;
                10'b0011101101: data = 24'b011100111011011001110001;
                10'b0011101110: data = 24'b011100111011011001110001;
                10'b0011101111: data = 24'b011100111011011001110001;
                10'b0011110000: data = 24'b011100111011011001110001;
                10'b0011110001: data = 24'b011100111011011001110001;
                10'b0011110010: data = 24'b011100111011011001110001;
                10'b0011110011: data = 24'b011100111011011001110001;
                10'b0011110100: data = 24'b011100111011011001110001;
                10'b0011110101: data = 24'b011100111011011001110001;
                10'b0011110110: data = 24'b011100111011011001110001;
                10'b0011110111: data = 24'b011100111011010001110001;
                10'b0011111000: data = 24'b011010111010000001101001;
                10'b0011111001: data = 24'b011010101001111001101000;
                10'b0011111010: data = 24'b011010101001111101101000;
                10'b0011111011: data = 24'b011010011001110101100111;
                10'b0011111100: data = 24'b010100100111100001010000;
                10'b0011111101: data = 24'b010011110111010101001110;
                10'b0011111110: data = 24'b010001000101101001000100;
                10'b0011111111: data = 24'b000000000000000000000000;
                10'b0100000000: data = 24'b000000000000000000000000;
                10'b0100000001: data = 24'b010001100101110001000101;
                10'b0100000010: data = 24'b010011110111010001001110;
                10'b0100000011: data = 24'b010100100111100001010000;
                10'b0100000100: data = 24'b011010011001110101100111;
                10'b0100000101: data = 24'b011010101001111101101000;
                10'b0100000110: data = 24'b011010101001110101101000;
                10'b0100000111: data = 24'b011011011010011101101011;
                10'b0100001000: data = 24'b011100111011011101110001;
                10'b0100001001: data = 24'b011100111011011001110001;
                10'b0100001010: data = 24'b011100111011011001110001;
                10'b0100001011: data = 24'b011100111011011001110001;
                10'b0100001100: data = 24'b011100111011011001110001;
                10'b0100001101: data = 24'b011100111011011001110001;
                10'b0100001110: data = 24'b011100111011011001110001;
                10'b0100001111: data = 24'b011100111011011001110001;
                10'b0100010000: data = 24'b011100111011011001110001;
                10'b0100010001: data = 24'b011100111011011001110001;
                10'b0100010010: data = 24'b011100111011011001110001;
                10'b0100010011: data = 24'b011100111011011001110001;
                10'b0100010100: data = 24'b011100111011011001110001;
                10'b0100010101: data = 24'b011100111011011001110001;
                10'b0100010110: data = 24'b011100111011011001110001;
                10'b0100010111: data = 24'b011100111011011001110001;
                10'b0100011000: data = 24'b011011001010010001101010;
                10'b0100011001: data = 24'b011010101001110101101000;
                10'b0100011010: data = 24'b011010101001111101101000;
                10'b0100011011: data = 24'b011010011001110101100111;
                10'b0100011100: data = 24'b010100100111100001010000;
                10'b0100011101: data = 24'b010011110111010001001110;
                10'b0100011110: data = 24'b010001100101110001000101;
                10'b0100011111: data = 24'b000000000000000000000000;
                10'b0100100000: data = 24'b000000000000000000000000;
                10'b0100100001: data = 24'b010000000101010001000000;
                10'b0100100010: data = 24'b010011110111010101001110;
                10'b0100100011: data = 24'b010100000111100001010000;
                10'b0100100100: data = 24'b011010011001110101100111;
                10'b0100100101: data = 24'b011010101001111101101000;
                10'b0100100110: data = 24'b011010011001110001100111;
                10'b0100100111: data = 24'b011011111010101001101101;
                10'b0100101000: data = 24'b011101001011100001110010;
                10'b0100101001: data = 24'b011100111011011001110001;
                10'b0100101010: data = 24'b011100111011011001110001;
                10'b0100101011: data = 24'b011100111011011001110001;
                10'b0100101100: data = 24'b011100111011011001110001;
                10'b0100101101: data = 24'b011100111011011001110001;
                10'b0100101110: data = 24'b011100111011011001110001;
                10'b0100101111: data = 24'b011100111011011001110001;
                10'b0100110000: data = 24'b011100111011011001110001;
                10'b0100110001: data = 24'b011100111011011001110001;
                10'b0100110010: data = 24'b011100111011011001110001;
                10'b0100110011: data = 24'b011100111011011001110001;
                10'b0100110100: data = 24'b011100111011011001110001;
                10'b0100110101: data = 24'b011100111011011001110001;
                10'b0100110110: data = 24'b011100111011011001110001;
                10'b0100110111: data = 24'b011101001011011101110010;
                10'b0100111000: data = 24'b011011101010100001101100;
                10'b0100111001: data = 24'b011010101001110101101000;
                10'b0100111010: data = 24'b011010101001111101101000;
                10'b0100111011: data = 24'b011010011001110101100111;
                10'b0100111100: data = 24'b010100000111100001010000;
                10'b0100111101: data = 24'b010011110111010101001110;
                10'b0100111110: data = 24'b010000000101010000111111;
                10'b0100111111: data = 24'b000000000000000000000000;
                10'b0101000000: data = 24'b000000000000000000000000;
                10'b0101000001: data = 24'b001011100011111100101101;
                10'b0101000010: data = 24'b010100010111011101010000;
                10'b0101000011: data = 24'b010011100111010001001101;
                10'b0101000100: data = 24'b011010011001110001100111;
                10'b0101000101: data = 24'b011010111001111101101001;
                10'b0101000110: data = 24'b011010011001110001100111;
                10'b0101000111: data = 24'b011011111010100101101101;
                10'b0101001000: data = 24'b011101001011100001110010;
                10'b0101001001: data = 24'b011100111011011001110001;
                10'b0101001010: data = 24'b011100111011011001110001;
                10'b0101001011: data = 24'b011100111011011001110001;
                10'b0101001100: data = 24'b011100111011011001110001;
                10'b0101001101: data = 24'b011100111011011001110001;
                10'b0101001110: data = 24'b011100111011011001110001;
                10'b0101001111: data = 24'b011100111011011001110001;
                10'b0101010000: data = 24'b011100111011011001110001;
                10'b0101010001: data = 24'b011100111011011001110001;
                10'b0101010010: data = 24'b011100111011011001110001;
                10'b0101010011: data = 24'b011100111011011001110001;
                10'b0101010100: data = 24'b011100111011011001110001;
                10'b0101010101: data = 24'b011100111011011001110001;
                10'b0101010110: data = 24'b011100111011011001110001;
                10'b0101010111: data = 24'b011101001011100001110010;
                10'b0101011000: data = 24'b011011111010101001101101;
                10'b0101011001: data = 24'b011010011001110001100111;
                10'b0101011010: data = 24'b011010111001111101101001;
                10'b0101011011: data = 24'b011010011001110001100111;
                10'b0101011100: data = 24'b010011100111010001001101;
                10'b0101011101: data = 24'b010100010111011001010000;
                10'b0101011110: data = 24'b001011100011111100101101;
                10'b0101011111: data = 24'b000000000000000000000000;
                10'b0101100000: data = 24'b000000000000000000000000;
                10'b0101100001: data = 24'b001001100011100000100110;
                10'b0101100010: data = 24'b010100100111100001010001;
                10'b0101100011: data = 24'b010011010111000101001100;
                10'b0101100100: data = 24'b011001101001100001100100;
                10'b0101100101: data = 24'b011010111001111101101001;
                10'b0101100110: data = 24'b011010101001110101101000;
                10'b0101100111: data = 24'b011011001010010101101010;
                10'b0101101000: data = 24'b011100111011011001110001;
                10'b0101101001: data = 24'b011100111011011001110001;
                10'b0101101010: data = 24'b011100111011011001110001;
                10'b0101101011: data = 24'b011100111011011001110001;
                10'b0101101100: data = 24'b011100111011011001110001;
                10'b0101101101: data = 24'b011100111011011001110001;
                10'b0101101110: data = 24'b011100111011011001110001;
                10'b0101101111: data = 24'b011100111011011001110001;
                10'b0101110000: data = 24'b011100111011011001110001;
                10'b0101110001: data = 24'b011100111011011001110001;
                10'b0101110010: data = 24'b011100111011011001110001;
                10'b0101110011: data = 24'b011100111011011001110001;
                10'b0101110100: data = 24'b011100111011011001110001;
                10'b0101110101: data = 24'b011100111011011001110001;
                10'b0101110110: data = 24'b011100111011011001110001;
                10'b0101110111: data = 24'b011101001011011101110010;
                10'b0101111000: data = 24'b011011101010100001101100;
                10'b0101111001: data = 24'b011010011001110001100111;
                10'b0101111010: data = 24'b011010111001111101101001;
                10'b0101111011: data = 24'b011001101001100001100100;
                10'b0101111100: data = 24'b010011010111000101001100;
                10'b0101111101: data = 24'b010100100111100001010001;
                10'b0101111110: data = 24'b001001110011101000100111;
                10'b0101111111: data = 24'b000000000000000000000000;
                10'b0110000000: data = 24'b000000000000000000000000;
                10'b0110000001: data = 24'b001010000011010000101000;
                10'b0110000010: data = 24'b010100010111010101010000;
                10'b0110000011: data = 24'b010011010111000001001011;
                10'b0110000100: data = 24'b011000101001001001100000;
                10'b0110000101: data = 24'b011010111010000001101001;
                10'b0110000110: data = 24'b011010101001111001101000;
                10'b0110000111: data = 24'b011010111010000101101001;
                10'b0110001000: data = 24'b011100111011010101110001;
                10'b0110001001: data = 24'b011101001011100101110010;
                10'b0110001010: data = 24'b011101101011101101110011;
                10'b0110001011: data = 24'b011101011011101001110011;
                10'b0110001100: data = 24'b011100111011011001110001;
                10'b0110001101: data = 24'b011100111011011001110001;
                10'b0110001110: data = 24'b011100111011011001110001;
                10'b0110001111: data = 24'b011100111011011001110001;
                10'b0110010000: data = 24'b011100111011011001110001;
                10'b0110010001: data = 24'b011100111011011001110001;
                10'b0110010010: data = 24'b011100111011011001110001;
                10'b0110010011: data = 24'b011100111011011001110001;
                10'b0110010100: data = 24'b011101011011101001110011;
                10'b0110010101: data = 24'b011101101011101101110011;
                10'b0110010110: data = 24'b011101001011100001110010;
                10'b0110010111: data = 24'b011100111011011001110001;
                10'b0110011000: data = 24'b011011011010010001101011;
                10'b0110011001: data = 24'b011010101001110101101000;
                10'b0110011010: data = 24'b011010111010000001101001;
                10'b0110011011: data = 24'b011000101001001001100000;
                10'b0110011100: data = 24'b010011000111000001001011;
                10'b0110011101: data = 24'b010100110111011101010010;
                10'b0110011110: data = 24'b001011110011110100101110;
                10'b0110011111: data = 24'b000000000000000000000000;
                10'b0110100000: data = 24'b000000000000000000000000;
                10'b0110100001: data = 24'b000101000001011000010100;
                10'b0110100010: data = 24'b010011000110111001001011;
                10'b0110100011: data = 24'b010010110110111101001010;
                10'b0110100100: data = 24'b010111011000100101011011;
                10'b0110100101: data = 24'b011011001010000101101010;
                10'b0110100110: data = 24'b011010101001111001101000;
                10'b0110100111: data = 24'b011010101001111101101000;
                10'b0110101000: data = 24'b011100011011000001101111;
                10'b0110101001: data = 24'b011010101010100001101001;
                10'b0110101010: data = 24'b011000001001010101011110;
                10'b0110101011: data = 24'b011001001001101101100010;
                10'b0110101100: data = 24'b011100111011011001110001;
                10'b0110101101: data = 24'b011100111011011101110001;
                10'b0110101110: data = 24'b011100111011011001110001;
                10'b0110101111: data = 24'b011100111011011001110001;
                10'b0110110000: data = 24'b011100111011011001110001;
                10'b0110110001: data = 24'b011100111011011001110001;
                10'b0110110010: data = 24'b011100111011011101110001;
                10'b0110110011: data = 24'b011100111011011001110001;
                10'b0110110100: data = 24'b011001001001101101100010;
                10'b0110110101: data = 24'b011000001001010101011110;
                10'b0110110110: data = 24'b011010101010011101101001;
                10'b0110110111: data = 24'b011100101011001101110000;
                10'b0110111000: data = 24'b011010111010000001101001;
                10'b0110111001: data = 24'b011010101001111001101000;
                10'b0110111010: data = 24'b011011001010000101101010;
                10'b0110111011: data = 24'b010111011000100101011011;
                10'b0110111100: data = 24'b010010110110111101001010;
                10'b0110111101: data = 24'b010011010110111101001100;
                10'b0110111110: data = 24'b000101100001101000010110;
                10'b0110111111: data = 24'b000000000000000000000000;
                10'b0111000000: data = 24'b000000000000000000000000;
                10'b0111000001: data = 24'b000000110000010100000011;
                10'b0111000010: data = 24'b010010110110011101001010;
                10'b0111000011: data = 24'b010011010111000101001100;
                10'b0111000100: data = 24'b010101010111111001010100;
                10'b0111000101: data = 24'b011010111010000001101001;
                10'b0111000110: data = 24'b011010101001111001101000;
                10'b0111000111: data = 24'b011010111001111101101000;
                10'b0111001000: data = 24'b010110111000100001011001;
                10'b0111001001: data = 24'b010011110111010001001110;
                10'b0111001010: data = 24'b010100100111010001010001;
                10'b0111001011: data = 24'b010011010110111101001100;
                10'b0111001100: data = 24'b011000101001100001100000;
                10'b0111001101: data = 24'b011101011011100101110011;
                10'b0111001110: data = 24'b011100111011011001110001;
                10'b0111001111: data = 24'b011100111011011001110001;
                10'b0111010000: data = 24'b011100111011011001110001;
                10'b0111010001: data = 24'b011100111011011001110001;
                10'b0111010010: data = 24'b011101011011100101110011;
                10'b0111010011: data = 24'b011000101001100001100000;
                10'b0111010100: data = 24'b010011010110111101001100;
                10'b0111010101: data = 24'b010100100111010001010001;
                10'b0111010110: data = 24'b010011110111001101001110;
                10'b0111010111: data = 24'b010110111000100101011010;
                10'b0111011000: data = 24'b011010111001111101101000;
                10'b0111011001: data = 24'b011010101001111001101000;
                10'b0111011010: data = 24'b011010111010000001101001;
                10'b0111011011: data = 24'b010101010111111001010100;
                10'b0111011100: data = 24'b010011000111000001001011;
                10'b0111011101: data = 24'b010011100110110101001101;
                10'b0111011110: data = 24'b000001000000010100000100;
                10'b0111011111: data = 24'b000000000000000000000000;
                10'b0111100000: data = 24'b000000000000000000000000;
                10'b0111100001: data = 24'b000000100000001000000010;
                10'b0111100010: data = 24'b001101110100101000110111;
                10'b0111100011: data = 24'b010100010111011101010000;
                10'b0111100100: data = 24'b010011100111001101001101;
                10'b0111100101: data = 24'b011001111001100101100101;
                10'b0111100110: data = 24'b011011001010000101101010;
                10'b0111100111: data = 24'b011000011001000101100000;
                10'b0111101000: data = 24'b010011110111001101001111;
                10'b0111101001: data = 24'b010111000111111101011011;
                10'b0111101010: data = 24'b011000001000001001011111;
                10'b0111101011: data = 24'b010110010111101101011000;
                10'b0111101100: data = 24'b010100010111101001010000;
                10'b0111101101: data = 24'b011100101011010001110000;
                10'b0111101110: data = 24'b011100111011011101110001;
                10'b0111101111: data = 24'b011100111011011001110001;
                10'b0111110000: data = 24'b011100111011011001110001;
                10'b0111110001: data = 24'b011100111011011101110001;
                10'b0111110010: data = 24'b011100101011010001110000;
                10'b0111110011: data = 24'b010100100111101001010001;
                10'b0111110100: data = 24'b010110010111101101011000;
                10'b0111110101: data = 24'b011000001000001001011111;
                10'b0111110110: data = 24'b010111000111111101011011;
                10'b0111110111: data = 24'b010011110111001001001111;
                10'b0111111000: data = 24'b011000011001000101100000;
                10'b0111111001: data = 24'b011011001010000101101010;
                10'b0111111010: data = 24'b011001111001100101100101;
                10'b0111111011: data = 24'b010011100111001101001101;
                10'b0111111100: data = 24'b010100000111011101001111;
                10'b0111111101: data = 24'b001110110100111100111010;
                10'b0111111110: data = 24'b000000100000001000000010;
                10'b0111111111: data = 24'b000000000000000000000000;
                10'b1000000000: data = 24'b000000000000000000000000;
                10'b1000000001: data = 24'b000000000000000000000000;
                10'b1000000010: data = 24'b001001100011000000100110;
                10'b1000000011: data = 24'b010100000111010001001111;
                10'b1000000100: data = 24'b010010110110111001001010;
                10'b1000000101: data = 24'b010111011000101101011100;
                10'b1000000110: data = 24'b011011101010010001101100;
                10'b1000000111: data = 24'b010110111000011101011001;
                10'b1000001000: data = 24'b010100110111010101010010;
                10'b1000001001: data = 24'b011000011000010001100000;
                10'b1000001010: data = 24'b011000011000010101100000;
                10'b1000001011: data = 24'b010111111000001001011110;
                10'b1000001100: data = 24'b010011110111010001001111;
                10'b1000001101: data = 24'b011010111010100001101001;
                10'b1000001110: data = 24'b011101011011100001110010;
                10'b1000001111: data = 24'b011100111011011001110001;
                10'b1000010000: data = 24'b011100111011011001110001;
                10'b1000010001: data = 24'b011101011011100001110010;
                10'b1000010010: data = 24'b011010111010100001101001;
                10'b1000010011: data = 24'b010011110111010001001111;
                10'b1000010100: data = 24'b010111111000001001011110;
                10'b1000010101: data = 24'b011000011000010101100000;
                10'b1000010110: data = 24'b011000011000010001100000;
                10'b1000010111: data = 24'b010100110111010101010010;
                10'b1000011000: data = 24'b010110111000011101011001;
                10'b1000011001: data = 24'b011011101010010001101100;
                10'b1000011010: data = 24'b010111011000101101011100;
                10'b1000011011: data = 24'b010010110110111001001010;
                10'b1000011100: data = 24'b010100010111011001010000;
                10'b1000011101: data = 24'b001010010011010000101001;
                10'b1000011110: data = 24'b000000000000000000000000;
                10'b1000011111: data = 24'b000000000000000000000000;
                10'b1000100000: data = 24'b000000000000000000000000;
                10'b1000100001: data = 24'b000000000000000000000000;
                10'b1000100010: data = 24'b000010110000110000001010;
                10'b1000100011: data = 24'b010010010110100001001001;
                10'b1000100100: data = 24'b010011010111001001001100;
                10'b1000100101: data = 24'b010100100111100101010001;
                10'b1000100110: data = 24'b011011001010000101101010;
                10'b1000100111: data = 24'b010111001000100101011010;
                10'b1000101000: data = 24'b010100110111011001010010;
                10'b1000101001: data = 24'b010101110111011101010110;
                10'b1000101010: data = 24'b010010110110100001001010;
                10'b1000101011: data = 24'b010101100111011001010101;
                10'b1000101100: data = 24'b010100100111011001010010;
                10'b1000101101: data = 24'b011001001001110101100010;
                10'b1000101110: data = 24'b011101011011101001110011;
                10'b1000101111: data = 24'b011100111011011001110001;
                10'b1000110000: data = 24'b011100111011011001110001;
                10'b1000110001: data = 24'b011101011011101001110011;
                10'b1000110010: data = 24'b011001001001110101100010;
                10'b1000110011: data = 24'b010100100111011001010010;
                10'b1000110100: data = 24'b010101100111011001010101;
                10'b1000110101: data = 24'b010010110110100001001010;
                10'b1000110110: data = 24'b010101110111011101010110;
                10'b1000110111: data = 24'b010100110111011001010010;
                10'b1000111000: data = 24'b010111001000100101011010;
                10'b1000111001: data = 24'b011011001010000101101010;
                10'b1000111010: data = 24'b010100100111100101010001;
                10'b1000111011: data = 24'b010011010111000101001100;
                10'b1000111100: data = 24'b010011000110110001001011;
                10'b1000111101: data = 24'b000011000000111000001100;
                10'b1000111110: data = 24'b000000000000000000000000;
                10'b1000111111: data = 24'b000000000000000000000000;
                10'b1001000000: data = 24'b000000000000000000000000;
                10'b1001000001: data = 24'b000000010000000100000001;
                10'b1001000010: data = 24'b000000110000001100000011;
                10'b1001000011: data = 24'b001101100100011000110101;
                10'b1001000100: data = 24'b010100100111100001010001;
                10'b1001000101: data = 24'b010011000110111101001011;
                10'b1001000110: data = 24'b011000111001010001100001;
                10'b1001000111: data = 24'b011000101001001001100000;
                10'b1001001000: data = 24'b010010110110110001001010;
                10'b1001001001: data = 24'b001110100101000100111001;
                10'b1001001010: data = 24'b001100110100100100110010;
                10'b1001001011: data = 24'b001110100101000100111001;
                10'b1001001100: data = 24'b010010110110101001001010;
                10'b1001001101: data = 24'b011000011001011101100000;
                10'b1001001110: data = 24'b011101101011101101110100;
                10'b1001001111: data = 24'b011100111011011001110001;
                10'b1001010000: data = 24'b011100111011011001110001;
                10'b1001010001: data = 24'b011101101011101101110100;
                10'b1001010010: data = 24'b011000011001011101100000;
                10'b1001010011: data = 24'b010010110110101001001010;
                10'b1001010100: data = 24'b001110100101000100111001;
                10'b1001010101: data = 24'b001100110100100100110010;
                10'b1001010110: data = 24'b001110100101000100111001;
                10'b1001010111: data = 24'b010010110110110001001010;
                10'b1001011000: data = 24'b011000101001001001100000;
                10'b1001011001: data = 24'b011000111001010001100001;
                10'b1001011010: data = 24'b010011000110111101001011;
                10'b1001011011: data = 24'b010100100111100001010000;
                10'b1001011100: data = 24'b001110010100101000111001;
                10'b1001011101: data = 24'b000000110000001100000011;
                10'b1001011110: data = 24'b000000010000000100000001;
                10'b1001011111: data = 24'b000000000000000000000000;
                10'b1001100000: data = 24'b000000000000000000000000;
                10'b1001100001: data = 24'b000000010000000100000001;
                10'b1001100010: data = 24'b000000000000000000000000;
                10'b1001100011: data = 24'b000101100001100100010110;
                10'b1001100100: data = 24'b010011100110111101001101;
                10'b1001100101: data = 24'b010011000111000001001011;
                10'b1001100110: data = 24'b010101010111111001010011;
                10'b1001100111: data = 24'b011010001001101101100110;
                10'b1001101000: data = 24'b010000110110000101000010;
                10'b1001101001: data = 24'b001101010100101100110100;
                10'b1001101010: data = 24'b001101110100111000110110;
                10'b1001101011: data = 24'b001101010100101100110100;
                10'b1001101100: data = 24'b001111110101101100111110;
                10'b1001101101: data = 24'b011000011001010101100000;
                10'b1001101110: data = 24'b011101101011101101110100;
                10'b1001101111: data = 24'b011100111011011001110001;
                10'b1001110000: data = 24'b011100111011011001110001;
                10'b1001110001: data = 24'b011101101011101101110100;
                10'b1001110010: data = 24'b011000011001010101100000;
                10'b1001110011: data = 24'b001111110101101100111110;
                10'b1001110100: data = 24'b001101010100101100110100;
                10'b1001110101: data = 24'b001101110100111000110110;
                10'b1001110110: data = 24'b001101010100101100110100;
                10'b1001110111: data = 24'b010000110110000101000010;
                10'b1001111000: data = 24'b011010001001101101100110;
                10'b1001111001: data = 24'b010101010111111001010011;
                10'b1001111010: data = 24'b010010110110111101001010;
                10'b1001111011: data = 24'b010011110111001001001111;
                10'b1001111100: data = 24'b000110000001110100011000;
                10'b1001111101: data = 24'b000000000000000000000000;
                10'b1001111110: data = 24'b000000010000000100000001;
                10'b1001111111: data = 24'b000000000000000000000000;
                10'b1010000000: data = 24'b000000000000000000000000;
                10'b1010000001: data = 24'b000000010000000100000001;
                10'b1010000010: data = 24'b000000010000000100000001;
                10'b1010000011: data = 24'b000000100000001000000010;
                10'b1010000100: data = 24'b001110000100101000111000;
                10'b1010000101: data = 24'b010100100111100001010001;
                10'b1010000110: data = 24'b010010110110111101001011;
                10'b1010000111: data = 24'b011000101001001101100001;
                10'b1010001000: data = 24'b010011010111000101001100;
                10'b1010001001: data = 24'b001101000100100100110011;
                10'b1010001010: data = 24'b001101100100110100110101;
                10'b1010001011: data = 24'b001101100100101100110101;
                10'b1010001100: data = 24'b010000110110000101000010;
                10'b1010001101: data = 24'b011000011001011101100000;
                10'b1010001110: data = 24'b011101101011101101110100;
                10'b1010001111: data = 24'b011100111011011001110001;
                10'b1010010000: data = 24'b011100111011011001110001;
                10'b1010010001: data = 24'b011101101011101101110100;
                10'b1010010010: data = 24'b011000011001011001100000;
                10'b1010010011: data = 24'b010000110110000101000010;
                10'b1010010100: data = 24'b001101100100101100110101;
                10'b1010010101: data = 24'b001101100100110100110101;
                10'b1010010110: data = 24'b001101000100100100110011;
                10'b1010010111: data = 24'b010011100111000101001100;
                10'b1010011000: data = 24'b011000101001001101100001;
                10'b1010011001: data = 24'b010010110110111101001011;
                10'b1010011010: data = 24'b010100010111100001010000;
                10'b1010011011: data = 24'b001111000101000000111011;
                10'b1010011100: data = 24'b000000100000001000000010;
                10'b1010011101: data = 24'b000000010000000100000001;
                10'b1010011110: data = 24'b000000010000000100000001;
                10'b1010011111: data = 24'b000000000000000000000000;
                10'b1010100000: data = 24'b000000000000000000000000;
                10'b1010100001: data = 24'b000000010000000100000001;
                10'b1010100010: data = 24'b000000010000000100000001;
                10'b1010100011: data = 24'b000000000000000000000000;
                10'b1010100100: data = 24'b000101010001011100010101;
                10'b1010100101: data = 24'b010011010110110101001101;
                10'b1010100110: data = 24'b010011010111000101001100;
                10'b1010100111: data = 24'b010100110111101001010001;
                10'b1010101000: data = 24'b010111101000101101011100;
                10'b1010101001: data = 24'b001111100101100100111101;
                10'b1010101010: data = 24'b001110010101000000111000;
                10'b1010101011: data = 24'b010001110110001001000110;
                10'b1010101100: data = 24'b010100000111001001001111;
                10'b1010101101: data = 24'b011001011001110101100011;
                10'b1010101110: data = 24'b011101011011101001110011;
                10'b1010101111: data = 24'b011100111011011001110001;
                10'b1010110000: data = 24'b011100111011011001110001;
                10'b1010110001: data = 24'b011101011011101001110011;
                10'b1010110010: data = 24'b011001011001110101100011;
                10'b1010110011: data = 24'b010100000111001001001111;
                10'b1010110100: data = 24'b010001110110001001000110;
                10'b1010110101: data = 24'b001110010101000000111000;
                10'b1010110110: data = 24'b001111100101100100111101;
                10'b1010110111: data = 24'b010111101000110001011100;
                10'b1010111000: data = 24'b010100100111101001010010;
                10'b1010111001: data = 24'b010011010111000001001100;
                10'b1010111010: data = 24'b010011110111000001001110;
                10'b1010111011: data = 24'b000101100001101100010110;
                10'b1010111100: data = 24'b000000000000000000000000;
                10'b1010111101: data = 24'b000000010000000100000001;
                10'b1010111110: data = 24'b000000010000000100000001;
                10'b1010111111: data = 24'b000000000000000000000000;
                10'b1011000000: data = 24'b000000000000000000000000;
                10'b1011000001: data = 24'b000000010000000100000001;
                10'b1011000010: data = 24'b000000010000000100000001;
                10'b1011000011: data = 24'b000000010000000100000001;
                10'b1011000100: data = 24'b000000100000001000000010;
                10'b1011000101: data = 24'b001100110100001100110011;
                10'b1011000110: data = 24'b010100100111100001010001;
                10'b1011000111: data = 24'b010010110110111001001010;
                10'b1011001000: data = 24'b010111011000100101011011;
                10'b1011001001: data = 24'b010110111000100001011010;
                10'b1011001010: data = 24'b010011100111000101001101;
                10'b1011001011: data = 24'b010100100111010001010001;
                10'b1011001100: data = 24'b010101000111110101010011;
                10'b1011001101: data = 24'b011100001011000101101110;
                10'b1011001110: data = 24'b011101001011011101110010;
                10'b1011001111: data = 24'b011100111011011001110001;
                10'b1011010000: data = 24'b011100111011011001110001;
                10'b1011010001: data = 24'b011101001011011101110010;
                10'b1011010010: data = 24'b011100001011000101101110;
                10'b1011010011: data = 24'b010101000111110101010011;
                10'b1011010100: data = 24'b010100100111010001010001;
                10'b1011010101: data = 24'b010011100111000101001101;
                10'b1011010110: data = 24'b010110111000100001011010;
                10'b1011010111: data = 24'b010111011000100101011011;
                10'b1011011000: data = 24'b010010110110111001001010;
                10'b1011011001: data = 24'b010100100111100101010010;
                10'b1011011010: data = 24'b001101110100100000110110;
                10'b1011011011: data = 24'b000000100000001000000010;
                10'b1011011100: data = 24'b000000010000000100000001;
                10'b1011011101: data = 24'b000000010000000100000001;
                10'b1011011110: data = 24'b000000010000000100000001;
                10'b1011011111: data = 24'b000000000000000000000000;
                10'b1011100000: data = 24'b000000000000000000000000;
                10'b1011100001: data = 24'b000000000000000000000000;
                10'b1011100010: data = 24'b000000010000000100000001;
                10'b1011100011: data = 24'b000000010000000100000001;
                10'b1011100100: data = 24'b000000000000000000000000;
                10'b1011100101: data = 24'b000011000000110100001100;
                10'b1011100110: data = 24'b010010000110010001000111;
                10'b1011100111: data = 24'b010011110111010101001110;
                10'b1011101000: data = 24'b010011010111001001001100;
                10'b1011101001: data = 24'b011001011001011101100011;
                10'b1011101010: data = 24'b011000101001001101100001;
                10'b1011101011: data = 24'b010110111000011101011010;
                10'b1011101100: data = 24'b011010011010000001100111;
                10'b1011101101: data = 24'b011101011011100101110010;
                10'b1011101110: data = 24'b011100111011011001110001;
                10'b1011101111: data = 24'b011100111011011001110001;
                10'b1011110000: data = 24'b011100111011011001110001;
                10'b1011110001: data = 24'b011100111011011101110001;
                10'b1011110010: data = 24'b011100101011010001110000;
                10'b1011110011: data = 24'b011001111001101101100101;
                10'b1011110100: data = 24'b010110111000100001011010;
                10'b1011110101: data = 24'b011000101001001101100001;
                10'b1011110110: data = 24'b011001011001011101100011;
                10'b1011110111: data = 24'b010011010111001001001100;
                10'b1011111000: data = 24'b010011100111010001001101;
                10'b1011111001: data = 24'b010011000110100101001011;
                10'b1011111010: data = 24'b000011010000111000001101;
                10'b1011111011: data = 24'b000000000000000000000000;
                10'b1011111100: data = 24'b000000010000000100000001;
                10'b1011111101: data = 24'b000000010000000100000001;
                10'b1011111110: data = 24'b000000010000000100000001;
                10'b1011111111: data = 24'b000000000000000000000000;
                10'b1100000000: data = 24'b000000000000000000000000;
                10'b1100000001: data = 24'b000000000000000000000000;
                10'b1100000010: data = 24'b000000000000000000000000;
                10'b1100000011: data = 24'b000000010000000100000001;
                10'b1100000100: data = 24'b000000010000000100000001;
                10'b1100000101: data = 24'b000000000000000000000000;
                10'b1100000110: data = 24'b001000100010101000100010;
                10'b1100000111: data = 24'b010100000111010001010000;
                10'b1100001000: data = 24'b010011000110111101001011;
                10'b1100001001: data = 24'b010100100111101001010001;
                10'b1100001010: data = 24'b011010101001111001101000;
                10'b1100001011: data = 24'b011011011010001001101011;
                10'b1100001100: data = 24'b011010111001111101101001;
                10'b1100001101: data = 24'b011011101010100101101100;
                10'b1100001110: data = 24'b011100111011011101110001;
                10'b1100001111: data = 24'b011100111011011101110001;
                10'b1100010000: data = 24'b011100111011011101110001;
                10'b1100010001: data = 24'b011100011011000101101111;
                10'b1100010010: data = 24'b011010111010000101101001;
                10'b1100010011: data = 24'b011010101001111001101000;
                10'b1100010100: data = 24'b011011011010001001101011;
                10'b1100010101: data = 24'b011010101001111001101000;
                10'b1100010110: data = 24'b010100100111101001010001;
                10'b1100010111: data = 24'b010010110110111101001010;
                10'b1100011000: data = 24'b010100100111011001010001;
                10'b1100011001: data = 24'b001001010010111000100101;
                10'b1100011010: data = 24'b000000000000000000000000;
                10'b1100011011: data = 24'b000000010000000100000001;
                10'b1100011100: data = 24'b000000000000000000000000;
                10'b1100011101: data = 24'b000000000000000000000000;
                10'b1100011110: data = 24'b000000000000000000000000;
                10'b1100011111: data = 24'b000000000000000000000000;
                10'b1100100000: data = 24'b000000000000000000000000;
                10'b1100100001: data = 24'b000000000000000000000000;
                10'b1100100010: data = 24'b000000000000000000000000;
                10'b1100100011: data = 24'b000000010000000100000001;
                10'b1100100100: data = 24'b000000010000000100000001;
                10'b1100100101: data = 24'b000000010000000100000001;
                10'b1100100110: data = 24'b000001010000010100000101;
                10'b1100100111: data = 24'b001110000100100100111000;
                10'b1100101000: data = 24'b010100110111101001010010;
                10'b1100101001: data = 24'b010010100110111001001001;
                10'b1100101010: data = 24'b010101100111111101010100;
                10'b1100101011: data = 24'b011010101001111101101001;
                10'b1100101100: data = 24'b011010111001111101101001;
                10'b1100101101: data = 24'b011010101001110101101000;
                10'b1100101110: data = 24'b011001111001011101100101;
                10'b1100101111: data = 24'b011011001010001001101010;
                10'b1100110000: data = 24'b011010111010000001101001;
                10'b1100110001: data = 24'b011001101001010001100100;
                10'b1100110010: data = 24'b011010101001110101101000;
                10'b1100110011: data = 24'b011010111001111101101001;
                10'b1100110100: data = 24'b011010101001111101101001;
                10'b1100110101: data = 24'b010101100111111101010100;
                10'b1100110110: data = 24'b010010100110111001001001;
                10'b1100110111: data = 24'b010100110111101001010010;
                10'b1100111000: data = 24'b001111010101000000111101;
                10'b1100111001: data = 24'b000001010000010100000101;
                10'b1100111010: data = 24'b000000010000000100000001;
                10'b1100111011: data = 24'b000000010000000100000001;
                10'b1100111100: data = 24'b000000000000000000000000;
                10'b1100111101: data = 24'b000000000000000000000000;
                10'b1100111110: data = 24'b000000000000000000000000;
                10'b1100111111: data = 24'b000000000000000000000000;
                10'b1101000000: data = 24'b000000000000000000000000;
                10'b1101000001: data = 24'b000000000000000000000000;
                10'b1101000010: data = 24'b000000000000000000000000;
                10'b1101000011: data = 24'b000000000000000000000000;
                10'b1101000100: data = 24'b000000010000000100000001;
                10'b1101000101: data = 24'b000000010000000100000001;
                10'b1101000110: data = 24'b000000000000000000000000;
                10'b1101000111: data = 24'b000010100000101100001001;
                10'b1101001000: data = 24'b010000110101110001000011;
                10'b1101001001: data = 24'b010100010111100001010000;
                10'b1101001010: data = 24'b010010100110110101001001;
                10'b1101001011: data = 24'b010110001000000101010110;
                10'b1101001100: data = 24'b011010111001111101101001;
                10'b1101001101: data = 24'b011010111001111001101001;
                10'b1101001110: data = 24'b010111011000000001011100;
                10'b1101001111: data = 24'b011001001001000001100010;
                10'b1101010000: data = 24'b011001001001000101100010;
                10'b1101010001: data = 24'b010111011000000001011101;
                10'b1101010010: data = 24'b011010111001111001101001;
                10'b1101010011: data = 24'b011010111001111101101001;
                10'b1101010100: data = 24'b010110001000000101010110;
                10'b1101010101: data = 24'b010010100110110101001001;
                10'b1101010110: data = 24'b010100010111011101010000;
                10'b1101010111: data = 24'b010001010101111101000101;
                10'b1101011000: data = 24'b000010100000110000001010;
                10'b1101011001: data = 24'b000000000000000000000000;
                10'b1101011010: data = 24'b000000010000000100000001;
                10'b1101011011: data = 24'b000000000000000000000000;
                10'b1101011100: data = 24'b000000000000000000000000;
                10'b1101011101: data = 24'b000000000000000000000000;
                10'b1101011110: data = 24'b000000000000000000000000;
                10'b1101011111: data = 24'b000000000000000000000000;
                10'b1101100000: data = 24'b000000000000000000000000;
                10'b1101100001: data = 24'b000000000000000000000000;
                10'b1101100010: data = 24'b000000000000000000000000;
                10'b1101100011: data = 24'b000000000000000000000000;
                10'b1101100100: data = 24'b000000000000000000000000;
                10'b1101100101: data = 24'b000000010000000100000001;
                10'b1101100110: data = 24'b000000010000000100000001;
                10'b1101100111: data = 24'b000000000000000000000000;
                10'b1101101000: data = 24'b000101100001100000010110;
                10'b1101101001: data = 24'b010010100110010001001010;
                10'b1101101010: data = 24'b010100010111011101010000;
                10'b1101101011: data = 24'b010010110110111001001010;
                10'b1101101100: data = 24'b010101010111110101010011;
                10'b1101101101: data = 24'b011001011001011001100011;
                10'b1101101110: data = 24'b011001111001011001100101;
                10'b1101101111: data = 24'b011010101001110101101000;
                10'b1101110000: data = 24'b011010101001110101101000;
                10'b1101110001: data = 24'b011001111001011001100101;
                10'b1101110010: data = 24'b011001011001011001100011;
                10'b1101110011: data = 24'b010101010111110101010011;
                10'b1101110100: data = 24'b010010110110111001001010;
                10'b1101110101: data = 24'b010100010111011001010000;
                10'b1101110110: data = 24'b010011100110101101001101;
                10'b1101110111: data = 24'b000110010001101100011001;
                10'b1101111000: data = 24'b000000000000000000000000;
                10'b1101111001: data = 24'b000000010000000100000001;
                10'b1101111010: data = 24'b000000010000000100000001;
                10'b1101111011: data = 24'b000000000000000000000000;
                10'b1101111100: data = 24'b000000000000000000000000;
                10'b1101111101: data = 24'b000000000000000000000000;
                10'b1101111110: data = 24'b000000000000000000000000;
                10'b1101111111: data = 24'b000000000000000000000000;
                10'b1110000000: data = 24'b000000000000000000000000;
                10'b1110000001: data = 24'b000000000000000000000000;
                10'b1110000010: data = 24'b000000000000000000000000;
                10'b1110000011: data = 24'b000000000000000000000000;
                10'b1110000100: data = 24'b000000000000000000000000;
                10'b1110000101: data = 24'b000000010000000100000001;
                10'b1110000110: data = 24'b000000010000000100000001;
                10'b1110000111: data = 24'b000000010000000100000001;
                10'b1110001000: data = 24'b000000000000000000000000;
                10'b1110001001: data = 24'b000110010001110100011001;
                10'b1110001010: data = 24'b010010100110010001001001;
                10'b1110001011: data = 24'b010100100111100001010001;
                10'b1110001100: data = 24'b010010110110111101001010;
                10'b1110001101: data = 24'b010011010111001001001100;
                10'b1110001110: data = 24'b010101111000000101010101;
                10'b1110001111: data = 24'b010110111000100001011010;
                10'b1110010000: data = 24'b010110111000100001011010;
                10'b1110010001: data = 24'b010101111000000101010101;
                10'b1110010010: data = 24'b010011010111001001001100;
                10'b1110010011: data = 24'b010010110110111001001010;
                10'b1110010100: data = 24'b010100010111100001010000;
                10'b1110010101: data = 24'b010011010110100101001100;
                10'b1110010110: data = 24'b000111010010001100011101;
                10'b1110010111: data = 24'b000000000000000000000000;
                10'b1110011000: data = 24'b000000010000000100000001;
                10'b1110011001: data = 24'b000000000000000000000000;
                10'b1110011010: data = 24'b000000000000000000000000;
                10'b1110011011: data = 24'b000000000000000000000000;
                10'b1110011100: data = 24'b000000000000000000000000;
                10'b1110011101: data = 24'b000000000000000000000000;
                10'b1110011110: data = 24'b000000000000000000000000;
                10'b1110011111: data = 24'b000000000000000000000000;
                10'b1110100000: data = 24'b000000000000000000000000;
                10'b1110100001: data = 24'b000000000000000000000000;
                10'b1110100010: data = 24'b000000000000000000000000;
                10'b1110100011: data = 24'b000000000000000000000000;
                10'b1110100100: data = 24'b000000000000000000000000;
                10'b1110100101: data = 24'b000000000000000000000000;
                10'b1110100110: data = 24'b000000000000000000000000;
                10'b1110100111: data = 24'b000000010000000100000001;
                10'b1110101000: data = 24'b000000010000000100000001;
                10'b1110101001: data = 24'b000000000000000000000000;
                10'b1110101010: data = 24'b000100110001010100010011;
                10'b1110101011: data = 24'b010000000101010100111111;
                10'b1110101100: data = 24'b010100100111011001010001;
                10'b1110101101: data = 24'b010100000111011001001111;
                10'b1110101110: data = 24'b010011000110111101001011;
                10'b1110101111: data = 24'b010010110110111101001010;
                10'b1110110000: data = 24'b010010110110111101001010;
                10'b1110110001: data = 24'b010011000110111101001011;
                10'b1110110010: data = 24'b010100000111011001001111;
                10'b1110110011: data = 24'b010100110111100001010010;
                10'b1110110100: data = 24'b010000100101101101000010;
                10'b1110110101: data = 24'b000101100001100000010101;
                10'b1110110110: data = 24'b000000000000000000000000;
                10'b1110110111: data = 24'b000000010000000100000001;
                10'b1110111000: data = 24'b000000010000000100000001;
                10'b1110111001: data = 24'b000000000000000000000000;
                10'b1110111010: data = 24'b000000000000000000000000;
                10'b1110111011: data = 24'b000000000000000000000000;
                10'b1110111100: data = 24'b000000000000000000000000;
                10'b1110111101: data = 24'b000000000000000000000000;
                10'b1110111110: data = 24'b000000000000000000000000;
                10'b1110111111: data = 24'b000000000000000000000000;
                10'b1111000000: data = 24'b000000000000000000000000;
                10'b1111000001: data = 24'b000000010000000100000001;
                10'b1111000010: data = 24'b000000000000000000000000;
                10'b1111000011: data = 24'b000000000000000000000000;
                10'b1111000100: data = 24'b000000000000000000000000;
                10'b1111000101: data = 24'b000000000000000000000000;
                10'b1111000110: data = 24'b000000000000000000000000;
                10'b1111000111: data = 24'b000000010000000100000001;
                10'b1111001000: data = 24'b000000010000000100000001;
                10'b1111001001: data = 24'b000000010000000100000001;
                10'b1111001010: data = 24'b000000000000000000000000;
                10'b1111001011: data = 24'b000000010000000100000001;
                10'b1111001100: data = 24'b000111100010100000011110;
                10'b1111001101: data = 24'b010000000101011100111111;
                10'b1111001110: data = 24'b010010110110110101001010;
                10'b1111001111: data = 24'b010010000110101001000111;
                10'b1111010000: data = 24'b010010000110101001000111;
                10'b1111010001: data = 24'b010010110110110101001010;
                10'b1111010010: data = 24'b010000000101011100111111;
                10'b1111010011: data = 24'b001000110010110100100010;
                10'b1111010100: data = 24'b000000010000000100000001;
                10'b1111010101: data = 24'b000000000000000000000000;
                10'b1111010110: data = 24'b000000010000000100000001;
                10'b1111010111: data = 24'b000000010000000100000001;
                10'b1111011000: data = 24'b000000010000000100000001;
                10'b1111011001: data = 24'b000000000000000000000000;
                10'b1111011010: data = 24'b000000000000000000000000;
                10'b1111011011: data = 24'b000000000000000000000000;
                10'b1111011100: data = 24'b000000000000000000000000;
                10'b1111011101: data = 24'b000000000000000000000000;
                10'b1111011110: data = 24'b000000000000000000000000;
                10'b1111011111: data = 24'b000000000000000000000000;
                10'b1111100000: data = 24'b000000000000000000000000;
                10'b1111100001: data = 24'b000000000000000000000000;
                10'b1111100010: data = 24'b000000000000000000000000;
                10'b1111100011: data = 24'b000000000000000000000000;
                10'b1111100100: data = 24'b000000000000000000000000;
                10'b1111100101: data = 24'b000000000000000000000000;
                10'b1111100110: data = 24'b000000000000000000000000;
                10'b1111100111: data = 24'b000000000000000000000000;
                10'b1111101000: data = 24'b000000000000000000000000;
                10'b1111101001: data = 24'b000000000000000000000000;
                10'b1111101010: data = 24'b000000000000000000000000;
                10'b1111101011: data = 24'b000000000000000000000000;
                10'b1111101100: data = 24'b000000000000000000000000;
                10'b1111101101: data = 24'b000000000000000000000000;
                10'b1111101110: data = 24'b000000000000000000000000;
                10'b1111101111: data = 24'b000000000000000000000000;
                10'b1111110000: data = 24'b000000000000000000000000;
                10'b1111110001: data = 24'b000000000000000000000000;
                10'b1111110010: data = 24'b000000000000000000000000;
                10'b1111110011: data = 24'b000000000000000000000000;
                10'b1111110100: data = 24'b000000000000000000000000;
                10'b1111110101: data = 24'b000000000000000000000000;
                10'b1111110110: data = 24'b000000000000000000000000;
                10'b1111110111: data = 24'b000000000000000000000000;
                10'b1111111000: data = 24'b000000000000000000000000;
                10'b1111111001: data = 24'b000000000000000000000000;
                10'b1111111010: data = 24'b000000000000000000000000;
                10'b1111111011: data = 24'b000000000000000000000000;
                10'b1111111100: data = 24'b000000000000000000000000;
                10'b1111111101: data = 24'b000000000000000000000000;
                10'b1111111110: data = 24'b000000000000000000000000;
                10'b1111111111: data = 24'b000000000000000000000000;
        endcase
        end
endmodule